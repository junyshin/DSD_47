entity g47_testbed is
  port (
  clock
  ) ;
end entity ; -- g47_testbed

architecture arch of g47_testbed is



begin



end architecture ; -- arch
