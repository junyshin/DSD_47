library ieee;
use ieee.std_logic_1164.all;

entity g47_enigma is
  port (
    clock
  ) ;
end entity ; -- g47_enigma

architecture arch of g47_enigma is

begin

end architecture ; -- arch
